// ---------------------- Full Adder de 1 bit ----------------------
module full_adder_1_bit (
    input  logic A,       // Entrada A
    input  logic B,       // Entrada B
    input  logic Cin,     // Acarreo de entrada
    output logic Sum,     // Suma
    output logic Cout     // Acarreo de salida
);

    // Resultado de la suma
    assign Sum  = A ^ B ^ Cin;     
	// Resultado de la suma	 (Acarreo de salida)
    assign Cout = (A & B) | (Cin & (A ^ B)); 

endmodule